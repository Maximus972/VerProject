module neg(
    input a,
    output c
);

    assign c = ~a;

endmodule;